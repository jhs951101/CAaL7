
module AdderLogic(ac_data, inp_r, dr_data, out);

input [15:0] ac_data;
input [7:0] inp_r;
input [15:0] dr_data;
output [15:0] out;
reg [15:0] out;

endmodule
