
module EFlipFlop(eff_in);

input eff_in;

reg eff_r;



endmodule
